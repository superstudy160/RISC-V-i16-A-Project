parameter MultiplicationOverflowIdx = 0;
parameter DivisionHasRemainderIdx = 1;
parameter DivisionByZeroIdx = 2;
parameter NoFlagsIdx = 3;