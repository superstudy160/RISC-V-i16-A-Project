module multiplication (
    input [0:15] M1,
    input [0:15] M2
);
    
endmodule