module ALU #(parameter l=16) (
	input [lv:0] A,
	input [lv:0] B,
	input [2:0] Operation,
	output [lv:0] R,
)

parameter lv = l-1;

// TODO: implement ALU

endmodule //ALU