module multiplication (
    
);
    
endmodule