module RISCV(
    input clk
);
    
endmodule //RISCV
