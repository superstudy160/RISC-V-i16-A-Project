module B(
	input a, 
	output wire b
);

	assign b = ~a;

endmodule