module Division #(parameter l=16) (
    input [lv:0] A,
    input [lv:0] B,
    output [lv:0] Quotient,
    output [lv:0] Remainder,
    output reg DivByZero
);

parameter lv = l-1;

// TODO: Implement the division
    
endmodule //Division
